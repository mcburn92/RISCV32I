module alu_tb ();
reg [31:0] opA, opB;
reg clk;
reg [3:0] aluOp;
wire[31:0] out;

alu steve (opA, opB, aluOp, clk, out);

initial begin
clk <=0;
opA<= 32'd15;
opB<= 32'd2;
aluOp<=4'b0000;
end

always #5 clk=~clk;

initial begin
#10
#10
aluOp<=4'b1000;
#10
aluOp<=4'b0111;
#10
aluOp<=4'b0110;
#10
aluOp<=4'b0100;
#10
aluOp<=4'b0001;
#10
aluOp<=4'b0101;
#10 $stop;
end

endmodule
